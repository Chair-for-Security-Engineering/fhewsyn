// Copyright 2021 Google LLC
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
module ReverseString(
  input wire [63:0] my_string,
  output wire [63:0] out
);
  wire [7:0] my_string_unflattened[0:7];
  assign my_string_unflattened[0] = my_string[7:0];
  assign my_string_unflattened[1] = my_string[15:8];
  assign my_string_unflattened[2] = my_string[23:16];
  assign my_string_unflattened[3] = my_string[31:24];
  assign my_string_unflattened[4] = my_string[39:32];
  assign my_string_unflattened[5] = my_string[47:40];
  assign my_string_unflattened[6] = my_string[55:48];
  assign my_string_unflattened[7] = my_string[63:56];
  wire [7:0] array_index_1736;
  wire [7:0] array_index_1740;
  wire [7:0] array_index_1747;
  wire [7:0] array_index_1754;
  wire [7:0] array_index_1761;
  wire [7:0] array_index_1767;
  wire [7:0] array_index_1779;
  wire [31:0] and_1790;
  wire [31:0] add_1792;
  wire [30:0] add_1797;
  wire [7:0] array_update_1799[0:7];
  wire [31:0] concat_1802;
  wire [7:0] array_update_1803[0:7];
  wire sgt_1804;
  wire [7:0] sel_1809[0:7];
  wire [31:0] add_1813;
  wire [7:0] array_update_1814[0:7];
  wire [7:0] array_update_1821[0:7];
  wire [29:0] add_1823;
  wire sgt_1825;
  wire [31:0] concat_1830;
  wire [7:0] sel_1831[0:7];
  wire [7:0] array_update_1838[0:7];
  wire [7:0] array_update_1845[0:7];
  wire [31:0] add_1848;
  wire sgt_1849;
  wire [7:0] sel_1858[0:7];
  wire [30:0] add_1864;
  wire [7:0] array_update_1867[0:7];
  wire [31:0] concat_1871;
  wire [7:0] array_update_1875[0:7];
  wire sgt_1881;
  wire [7:0] sel_1891[0:7];
  wire [31:0] add_1898;
  wire [7:0] array_update_1901[0:7];
  wire [7:0] array_update_1911[0:7];
  wire sgt_1918;
  wire [7:0] sel_1928[0:7];
  wire [7:0] array_update_1938[0:7];
  wire [7:0] array_update_1946[0:7];
  wire sgt_1950;
  wire [7:0] sel_1956[0:7];
  wire [7:0] array_update_1962[0:7];
  wire [7:0] array_update_1965[0:7];
  wire [7:0] sel_1966[0:7];
  assign array_index_1736 = my_string_unflattened[3'h6];
  assign array_index_1740 = my_string_unflattened[3'h5];
  assign array_index_1747 = my_string_unflattened[3'h4];
  assign array_index_1754 = my_string_unflattened[3'h3];
  assign array_index_1761 = my_string_unflattened[3'h2];
  assign array_index_1767 = my_string_unflattened[3'h1];
  assign array_index_1779 = my_string_unflattened[3'h0];
  assign and_1790 = {28'h000_0000, {{24{array_index_1767[7]}}, array_index_1767} == 32'h0000_0000 ? 4'h1 : ({{24{array_index_1761[7]}}, array_index_1761} == 32'h0000_0000 ? 4'h2 : ({{24{array_index_1754[7]}}, array_index_1754} == 32'h0000_0000 ? 4'h3 : ({{24{array_index_1747[7]}}, array_index_1747} == 32'h0000_0000 ? 4'h4 : ({{24{array_index_1740[7]}}, array_index_1740} == 32'h0000_0000 ? 4'h5 : ({{24{array_index_1736[7]}}, array_index_1736} == 32'h0000_0000 ? 4'h6 : ({{24{my_string_unflattened[3'h7][7]}}, my_string_unflattened[3'h7]} == 32'h0000_0000 ? 4'h7 : 4'h8))))))} & {32{{{24{array_index_1779[7]}}, array_index_1779} != 32'h0000_0000}};
  assign add_1792 = and_1790 + 32'hffff_ffff;
  assign add_1797 = and_1790[31:1] + 31'h7fff_ffff;
  assign array_update_1799[0] = my_string_unflattened[add_1792 > 32'h0000_0007 ? 32'h0000_0007 : add_1792];
  assign array_update_1799[1] = my_string_unflattened[1];
  assign array_update_1799[2] = my_string_unflattened[2];
  assign array_update_1799[3] = my_string_unflattened[3];
  assign array_update_1799[4] = my_string_unflattened[4];
  assign array_update_1799[5] = my_string_unflattened[5];
  assign array_update_1799[6] = my_string_unflattened[6];
  assign array_update_1799[7] = my_string_unflattened[7];
  assign concat_1802 = {add_1797, and_1790[0]};
  assign array_update_1803[0] = add_1792 == 32'h0000_0000 ? array_index_1779 : array_update_1799[0];
  assign array_update_1803[1] = add_1792 == 32'h0000_0001 ? array_index_1779 : array_update_1799[1];
  assign array_update_1803[2] = add_1792 == 32'h0000_0002 ? array_index_1779 : array_update_1799[2];
  assign array_update_1803[3] = add_1792 == 32'h0000_0003 ? array_index_1779 : array_update_1799[3];
  assign array_update_1803[4] = add_1792 == 32'h0000_0004 ? array_index_1779 : array_update_1799[4];
  assign array_update_1803[5] = add_1792 == 32'h0000_0005 ? array_index_1779 : array_update_1799[5];
  assign array_update_1803[6] = add_1792 == 32'h0000_0006 ? array_index_1779 : array_update_1799[6];
  assign array_update_1803[7] = add_1792 == 32'h0000_0007 ? array_index_1779 : array_update_1799[7];
  assign sgt_1804 = $signed(and_1790[4:1]) > $signed(4'h0);
  assign sel_1809[0] = sgt_1804 == 1'h0 ? my_string_unflattened[0] : array_update_1803[0];
  assign sel_1809[1] = sgt_1804 == 1'h0 ? my_string_unflattened[1] : array_update_1803[1];
  assign sel_1809[2] = sgt_1804 == 1'h0 ? my_string_unflattened[2] : array_update_1803[2];
  assign sel_1809[3] = sgt_1804 == 1'h0 ? my_string_unflattened[3] : array_update_1803[3];
  assign sel_1809[4] = sgt_1804 == 1'h0 ? my_string_unflattened[4] : array_update_1803[4];
  assign sel_1809[5] = sgt_1804 == 1'h0 ? my_string_unflattened[5] : array_update_1803[5];
  assign sel_1809[6] = sgt_1804 == 1'h0 ? my_string_unflattened[6] : array_update_1803[6];
  assign sel_1809[7] = sgt_1804 == 1'h0 ? my_string_unflattened[7] : array_update_1803[7];
  assign add_1813 = and_1790 + 32'hffff_fffd;
  assign array_update_1814[0] = sel_1809[0];
  assign array_update_1814[1] = sgt_1804 ? array_update_1803[concat_1802 > 32'h0000_0007 ? 32'h0000_0007 : concat_1802] : my_string_unflattened[concat_1802 > 32'h0000_0007 ? 32'h0000_0007 : concat_1802];
  assign array_update_1814[2] = sel_1809[2];
  assign array_update_1814[3] = sel_1809[3];
  assign array_update_1814[4] = sel_1809[4];
  assign array_update_1814[5] = sel_1809[5];
  assign array_update_1814[6] = sel_1809[6];
  assign array_update_1814[7] = sel_1809[7];
  assign array_update_1821[0] = concat_1802 == 32'h0000_0000 ? (sgt_1804 ? array_update_1803[3'h1] : array_index_1767) : array_update_1814[0];
  assign array_update_1821[1] = concat_1802 == 32'h0000_0001 ? (sgt_1804 ? array_update_1803[3'h1] : array_index_1767) : array_update_1814[1];
  assign array_update_1821[2] = concat_1802 == 32'h0000_0002 ? (sgt_1804 ? array_update_1803[3'h1] : array_index_1767) : array_update_1814[2];
  assign array_update_1821[3] = concat_1802 == 32'h0000_0003 ? (sgt_1804 ? array_update_1803[3'h1] : array_index_1767) : array_update_1814[3];
  assign array_update_1821[4] = concat_1802 == 32'h0000_0004 ? (sgt_1804 ? array_update_1803[3'h1] : array_index_1767) : array_update_1814[4];
  assign array_update_1821[5] = concat_1802 == 32'h0000_0005 ? (sgt_1804 ? array_update_1803[3'h1] : array_index_1767) : array_update_1814[5];
  assign array_update_1821[6] = concat_1802 == 32'h0000_0006 ? (sgt_1804 ? array_update_1803[3'h1] : array_index_1767) : array_update_1814[6];
  assign array_update_1821[7] = concat_1802 == 32'h0000_0007 ? (sgt_1804 ? array_update_1803[3'h1] : array_index_1767) : array_update_1814[7];
  assign add_1823 = and_1790[31:2] + 30'h3fff_ffff;
  assign sgt_1825 = $signed(and_1790[4:1]) > $signed(4'h1);
  assign concat_1830 = {add_1823, and_1790[1:0]};
  assign sel_1831[0] = sgt_1825 == 1'h0 ? sel_1809[0] : array_update_1821[0];
  assign sel_1831[1] = sgt_1825 == 1'h0 ? sel_1809[1] : array_update_1821[1];
  assign sel_1831[2] = sgt_1825 == 1'h0 ? sel_1809[2] : array_update_1821[2];
  assign sel_1831[3] = sgt_1825 == 1'h0 ? sel_1809[3] : array_update_1821[3];
  assign sel_1831[4] = sgt_1825 == 1'h0 ? sel_1809[4] : array_update_1821[4];
  assign sel_1831[5] = sgt_1825 == 1'h0 ? sel_1809[5] : array_update_1821[5];
  assign sel_1831[6] = sgt_1825 == 1'h0 ? sel_1809[6] : array_update_1821[6];
  assign sel_1831[7] = sgt_1825 == 1'h0 ? sel_1809[7] : array_update_1821[7];
  assign array_update_1838[0] = sel_1831[0];
  assign array_update_1838[1] = sel_1831[1];
  assign array_update_1838[2] = sgt_1825 ? array_update_1821[add_1813 > 32'h0000_0007 ? 32'h0000_0007 : add_1813] : (sgt_1804 ? array_update_1803[add_1813 > 32'h0000_0007 ? 32'h0000_0007 : add_1813] : my_string_unflattened[add_1813 > 32'h0000_0007 ? 32'h0000_0007 : add_1813]);
  assign array_update_1838[3] = sel_1831[3];
  assign array_update_1838[4] = sel_1831[4];
  assign array_update_1838[5] = sel_1831[5];
  assign array_update_1838[6] = sel_1831[6];
  assign array_update_1838[7] = sel_1831[7];
  assign array_update_1845[0] = add_1813 == 32'h0000_0000 ? (sgt_1825 ? array_update_1821[3'h2] : (sgt_1804 ? array_update_1803[3'h2] : array_index_1761)) : array_update_1838[0];
  assign array_update_1845[1] = add_1813 == 32'h0000_0001 ? (sgt_1825 ? array_update_1821[3'h2] : (sgt_1804 ? array_update_1803[3'h2] : array_index_1761)) : array_update_1838[1];
  assign array_update_1845[2] = add_1813 == 32'h0000_0002 ? (sgt_1825 ? array_update_1821[3'h2] : (sgt_1804 ? array_update_1803[3'h2] : array_index_1761)) : array_update_1838[2];
  assign array_update_1845[3] = add_1813 == 32'h0000_0003 ? (sgt_1825 ? array_update_1821[3'h2] : (sgt_1804 ? array_update_1803[3'h2] : array_index_1761)) : array_update_1838[3];
  assign array_update_1845[4] = add_1813 == 32'h0000_0004 ? (sgt_1825 ? array_update_1821[3'h2] : (sgt_1804 ? array_update_1803[3'h2] : array_index_1761)) : array_update_1838[4];
  assign array_update_1845[5] = add_1813 == 32'h0000_0005 ? (sgt_1825 ? array_update_1821[3'h2] : (sgt_1804 ? array_update_1803[3'h2] : array_index_1761)) : array_update_1838[5];
  assign array_update_1845[6] = add_1813 == 32'h0000_0006 ? (sgt_1825 ? array_update_1821[3'h2] : (sgt_1804 ? array_update_1803[3'h2] : array_index_1761)) : array_update_1838[6];
  assign array_update_1845[7] = add_1813 == 32'h0000_0007 ? (sgt_1825 ? array_update_1821[3'h2] : (sgt_1804 ? array_update_1803[3'h2] : array_index_1761)) : array_update_1838[7];
  assign add_1848 = and_1790 + 32'hffff_fffb;
  assign sgt_1849 = $signed(and_1790[4:1]) > $signed(4'h2);
  assign sel_1858[0] = sgt_1849 == 1'h0 ? sel_1831[0] : array_update_1845[0];
  assign sel_1858[1] = sgt_1849 == 1'h0 ? sel_1831[1] : array_update_1845[1];
  assign sel_1858[2] = sgt_1849 == 1'h0 ? sel_1831[2] : array_update_1845[2];
  assign sel_1858[3] = sgt_1849 == 1'h0 ? sel_1831[3] : array_update_1845[3];
  assign sel_1858[4] = sgt_1849 == 1'h0 ? sel_1831[4] : array_update_1845[4];
  assign sel_1858[5] = sgt_1849 == 1'h0 ? sel_1831[5] : array_update_1845[5];
  assign sel_1858[6] = sgt_1849 == 1'h0 ? sel_1831[6] : array_update_1845[6];
  assign sel_1858[7] = sgt_1849 == 1'h0 ? sel_1831[7] : array_update_1845[7];
  assign add_1864 = and_1790[31:1] + 31'h7fff_fffd;
  assign array_update_1867[0] = sel_1858[0];
  assign array_update_1867[1] = sel_1858[1];
  assign array_update_1867[2] = sel_1858[2];
  assign array_update_1867[3] = sgt_1849 ? array_update_1845[concat_1830 > 32'h0000_0007 ? 32'h0000_0007 : concat_1830] : (sgt_1825 ? array_update_1821[concat_1830 > 32'h0000_0007 ? 32'h0000_0007 : concat_1830] : (sgt_1804 ? array_update_1803[concat_1830 > 32'h0000_0007 ? 32'h0000_0007 : concat_1830] : my_string_unflattened[concat_1830 > 32'h0000_0007 ? 32'h0000_0007 : concat_1830]));
  assign array_update_1867[4] = sel_1858[4];
  assign array_update_1867[5] = sel_1858[5];
  assign array_update_1867[6] = sel_1858[6];
  assign array_update_1867[7] = sel_1858[7];
  assign concat_1871 = {add_1864, and_1790[0]};
  assign array_update_1875[0] = concat_1830 == 32'h0000_0000 ? (sgt_1849 ? array_update_1845[3'h3] : (sgt_1825 ? array_update_1821[3'h3] : (sgt_1804 ? array_update_1803[3'h3] : array_index_1754))) : array_update_1867[0];
  assign array_update_1875[1] = concat_1830 == 32'h0000_0001 ? (sgt_1849 ? array_update_1845[3'h3] : (sgt_1825 ? array_update_1821[3'h3] : (sgt_1804 ? array_update_1803[3'h3] : array_index_1754))) : array_update_1867[1];
  assign array_update_1875[2] = concat_1830 == 32'h0000_0002 ? (sgt_1849 ? array_update_1845[3'h3] : (sgt_1825 ? array_update_1821[3'h3] : (sgt_1804 ? array_update_1803[3'h3] : array_index_1754))) : array_update_1867[2];
  assign array_update_1875[3] = concat_1830 == 32'h0000_0003 ? (sgt_1849 ? array_update_1845[3'h3] : (sgt_1825 ? array_update_1821[3'h3] : (sgt_1804 ? array_update_1803[3'h3] : array_index_1754))) : array_update_1867[3];
  assign array_update_1875[4] = concat_1830 == 32'h0000_0004 ? (sgt_1849 ? array_update_1845[3'h3] : (sgt_1825 ? array_update_1821[3'h3] : (sgt_1804 ? array_update_1803[3'h3] : array_index_1754))) : array_update_1867[4];
  assign array_update_1875[5] = concat_1830 == 32'h0000_0005 ? (sgt_1849 ? array_update_1845[3'h3] : (sgt_1825 ? array_update_1821[3'h3] : (sgt_1804 ? array_update_1803[3'h3] : array_index_1754))) : array_update_1867[5];
  assign array_update_1875[6] = concat_1830 == 32'h0000_0006 ? (sgt_1849 ? array_update_1845[3'h3] : (sgt_1825 ? array_update_1821[3'h3] : (sgt_1804 ? array_update_1803[3'h3] : array_index_1754))) : array_update_1867[6];
  assign array_update_1875[7] = concat_1830 == 32'h0000_0007 ? (sgt_1849 ? array_update_1845[3'h3] : (sgt_1825 ? array_update_1821[3'h3] : (sgt_1804 ? array_update_1803[3'h3] : array_index_1754))) : array_update_1867[7];
  assign sgt_1881 = $signed(and_1790[4:1]) > $signed(4'h3);
  assign sel_1891[0] = sgt_1881 == 1'h0 ? sel_1858[0] : array_update_1875[0];
  assign sel_1891[1] = sgt_1881 == 1'h0 ? sel_1858[1] : array_update_1875[1];
  assign sel_1891[2] = sgt_1881 == 1'h0 ? sel_1858[2] : array_update_1875[2];
  assign sel_1891[3] = sgt_1881 == 1'h0 ? sel_1858[3] : array_update_1875[3];
  assign sel_1891[4] = sgt_1881 == 1'h0 ? sel_1858[4] : array_update_1875[4];
  assign sel_1891[5] = sgt_1881 == 1'h0 ? sel_1858[5] : array_update_1875[5];
  assign sel_1891[6] = sgt_1881 == 1'h0 ? sel_1858[6] : array_update_1875[6];
  assign sel_1891[7] = sgt_1881 == 1'h0 ? sel_1858[7] : array_update_1875[7];
  assign add_1898 = and_1790 + 32'hffff_fff9;
  assign array_update_1901[0] = sel_1891[0];
  assign array_update_1901[1] = sel_1891[1];
  assign array_update_1901[2] = sel_1891[2];
  assign array_update_1901[3] = sel_1891[3];
  assign array_update_1901[4] = sgt_1881 ? array_update_1875[add_1848 > 32'h0000_0007 ? 32'h0000_0007 : add_1848] : (sgt_1849 ? array_update_1845[add_1848 > 32'h0000_0007 ? 32'h0000_0007 : add_1848] : (sgt_1825 ? array_update_1821[add_1848 > 32'h0000_0007 ? 32'h0000_0007 : add_1848] : (sgt_1804 ? array_update_1803[add_1848 > 32'h0000_0007 ? 32'h0000_0007 : add_1848] : my_string_unflattened[add_1848 > 32'h0000_0007 ? 32'h0000_0007 : add_1848])));
  assign array_update_1901[5] = sel_1891[5];
  assign array_update_1901[6] = sel_1891[6];
  assign array_update_1901[7] = sel_1891[7];
  assign array_update_1911[0] = add_1848 == 32'h0000_0000 ? (sgt_1881 ? array_update_1875[3'h4] : (sgt_1849 ? array_update_1845[3'h4] : (sgt_1825 ? array_update_1821[3'h4] : (sgt_1804 ? array_update_1803[3'h4] : array_index_1747)))) : array_update_1901[0];
  assign array_update_1911[1] = add_1848 == 32'h0000_0001 ? (sgt_1881 ? array_update_1875[3'h4] : (sgt_1849 ? array_update_1845[3'h4] : (sgt_1825 ? array_update_1821[3'h4] : (sgt_1804 ? array_update_1803[3'h4] : array_index_1747)))) : array_update_1901[1];
  assign array_update_1911[2] = add_1848 == 32'h0000_0002 ? (sgt_1881 ? array_update_1875[3'h4] : (sgt_1849 ? array_update_1845[3'h4] : (sgt_1825 ? array_update_1821[3'h4] : (sgt_1804 ? array_update_1803[3'h4] : array_index_1747)))) : array_update_1901[2];
  assign array_update_1911[3] = add_1848 == 32'h0000_0003 ? (sgt_1881 ? array_update_1875[3'h4] : (sgt_1849 ? array_update_1845[3'h4] : (sgt_1825 ? array_update_1821[3'h4] : (sgt_1804 ? array_update_1803[3'h4] : array_index_1747)))) : array_update_1901[3];
  assign array_update_1911[4] = add_1848 == 32'h0000_0004 ? (sgt_1881 ? array_update_1875[3'h4] : (sgt_1849 ? array_update_1845[3'h4] : (sgt_1825 ? array_update_1821[3'h4] : (sgt_1804 ? array_update_1803[3'h4] : array_index_1747)))) : array_update_1901[4];
  assign array_update_1911[5] = add_1848 == 32'h0000_0005 ? (sgt_1881 ? array_update_1875[3'h4] : (sgt_1849 ? array_update_1845[3'h4] : (sgt_1825 ? array_update_1821[3'h4] : (sgt_1804 ? array_update_1803[3'h4] : array_index_1747)))) : array_update_1901[5];
  assign array_update_1911[6] = add_1848 == 32'h0000_0006 ? (sgt_1881 ? array_update_1875[3'h4] : (sgt_1849 ? array_update_1845[3'h4] : (sgt_1825 ? array_update_1821[3'h4] : (sgt_1804 ? array_update_1803[3'h4] : array_index_1747)))) : array_update_1901[6];
  assign array_update_1911[7] = add_1848 == 32'h0000_0007 ? (sgt_1881 ? array_update_1875[3'h4] : (sgt_1849 ? array_update_1845[3'h4] : (sgt_1825 ? array_update_1821[3'h4] : (sgt_1804 ? array_update_1803[3'h4] : array_index_1747)))) : array_update_1901[7];
  assign sgt_1918 = $signed(and_1790[4:1]) > $signed(4'h4);
  assign sel_1928[0] = sgt_1918 == 1'h0 ? sel_1891[0] : array_update_1911[0];
  assign sel_1928[1] = sgt_1918 == 1'h0 ? sel_1891[1] : array_update_1911[1];
  assign sel_1928[2] = sgt_1918 == 1'h0 ? sel_1891[2] : array_update_1911[2];
  assign sel_1928[3] = sgt_1918 == 1'h0 ? sel_1891[3] : array_update_1911[3];
  assign sel_1928[4] = sgt_1918 == 1'h0 ? sel_1891[4] : array_update_1911[4];
  assign sel_1928[5] = sgt_1918 == 1'h0 ? sel_1891[5] : array_update_1911[5];
  assign sel_1928[6] = sgt_1918 == 1'h0 ? sel_1891[6] : array_update_1911[6];
  assign sel_1928[7] = sgt_1918 == 1'h0 ? sel_1891[7] : array_update_1911[7];
  assign array_update_1938[0] = sel_1928[0];
  assign array_update_1938[1] = sel_1928[1];
  assign array_update_1938[2] = sel_1928[2];
  assign array_update_1938[3] = sel_1928[3];
  assign array_update_1938[4] = sel_1928[4];
  assign array_update_1938[5] = sgt_1918 ? array_update_1911[concat_1871 > 32'h0000_0007 ? 32'h0000_0007 : concat_1871] : (sgt_1881 ? array_update_1875[concat_1871 > 32'h0000_0007 ? 32'h0000_0007 : concat_1871] : (sgt_1849 ? array_update_1845[concat_1871 > 32'h0000_0007 ? 32'h0000_0007 : concat_1871] : (sgt_1825 ? array_update_1821[concat_1871 > 32'h0000_0007 ? 32'h0000_0007 : concat_1871] : (sgt_1804 ? array_update_1803[concat_1871 > 32'h0000_0007 ? 32'h0000_0007 : concat_1871] : my_string_unflattened[concat_1871 > 32'h0000_0007 ? 32'h0000_0007 : concat_1871]))));
  assign array_update_1938[6] = sel_1928[6];
  assign array_update_1938[7] = sel_1928[7];
  assign array_update_1946[0] = concat_1871 == 32'h0000_0000 ? (sgt_1918 ? array_update_1911[3'h5] : (sgt_1881 ? array_update_1875[3'h5] : (sgt_1849 ? array_update_1845[3'h5] : (sgt_1825 ? array_update_1821[3'h5] : (sgt_1804 ? array_update_1803[3'h5] : array_index_1740))))) : array_update_1938[0];
  assign array_update_1946[1] = concat_1871 == 32'h0000_0001 ? (sgt_1918 ? array_update_1911[3'h5] : (sgt_1881 ? array_update_1875[3'h5] : (sgt_1849 ? array_update_1845[3'h5] : (sgt_1825 ? array_update_1821[3'h5] : (sgt_1804 ? array_update_1803[3'h5] : array_index_1740))))) : array_update_1938[1];
  assign array_update_1946[2] = concat_1871 == 32'h0000_0002 ? (sgt_1918 ? array_update_1911[3'h5] : (sgt_1881 ? array_update_1875[3'h5] : (sgt_1849 ? array_update_1845[3'h5] : (sgt_1825 ? array_update_1821[3'h5] : (sgt_1804 ? array_update_1803[3'h5] : array_index_1740))))) : array_update_1938[2];
  assign array_update_1946[3] = concat_1871 == 32'h0000_0003 ? (sgt_1918 ? array_update_1911[3'h5] : (sgt_1881 ? array_update_1875[3'h5] : (sgt_1849 ? array_update_1845[3'h5] : (sgt_1825 ? array_update_1821[3'h5] : (sgt_1804 ? array_update_1803[3'h5] : array_index_1740))))) : array_update_1938[3];
  assign array_update_1946[4] = concat_1871 == 32'h0000_0004 ? (sgt_1918 ? array_update_1911[3'h5] : (sgt_1881 ? array_update_1875[3'h5] : (sgt_1849 ? array_update_1845[3'h5] : (sgt_1825 ? array_update_1821[3'h5] : (sgt_1804 ? array_update_1803[3'h5] : array_index_1740))))) : array_update_1938[4];
  assign array_update_1946[5] = concat_1871 == 32'h0000_0005 ? (sgt_1918 ? array_update_1911[3'h5] : (sgt_1881 ? array_update_1875[3'h5] : (sgt_1849 ? array_update_1845[3'h5] : (sgt_1825 ? array_update_1821[3'h5] : (sgt_1804 ? array_update_1803[3'h5] : array_index_1740))))) : array_update_1938[5];
  assign array_update_1946[6] = concat_1871 == 32'h0000_0006 ? (sgt_1918 ? array_update_1911[3'h5] : (sgt_1881 ? array_update_1875[3'h5] : (sgt_1849 ? array_update_1845[3'h5] : (sgt_1825 ? array_update_1821[3'h5] : (sgt_1804 ? array_update_1803[3'h5] : array_index_1740))))) : array_update_1938[6];
  assign array_update_1946[7] = concat_1871 == 32'h0000_0007 ? (sgt_1918 ? array_update_1911[3'h5] : (sgt_1881 ? array_update_1875[3'h5] : (sgt_1849 ? array_update_1845[3'h5] : (sgt_1825 ? array_update_1821[3'h5] : (sgt_1804 ? array_update_1803[3'h5] : array_index_1740))))) : array_update_1938[7];
  assign sgt_1950 = $signed(and_1790[4:1]) > $signed(4'h5);
  assign sel_1956[0] = sgt_1950 == 1'h0 ? sel_1928[0] : array_update_1946[0];
  assign sel_1956[1] = sgt_1950 == 1'h0 ? sel_1928[1] : array_update_1946[1];
  assign sel_1956[2] = sgt_1950 == 1'h0 ? sel_1928[2] : array_update_1946[2];
  assign sel_1956[3] = sgt_1950 == 1'h0 ? sel_1928[3] : array_update_1946[3];
  assign sel_1956[4] = sgt_1950 == 1'h0 ? sel_1928[4] : array_update_1946[4];
  assign sel_1956[5] = sgt_1950 == 1'h0 ? sel_1928[5] : array_update_1946[5];
  assign sel_1956[6] = sgt_1950 == 1'h0 ? sel_1928[6] : array_update_1946[6];
  assign sel_1956[7] = sgt_1950 == 1'h0 ? sel_1928[7] : array_update_1946[7];
  assign array_update_1962[0] = sel_1956[0];
  assign array_update_1962[1] = sel_1956[1];
  assign array_update_1962[2] = sel_1956[2];
  assign array_update_1962[3] = sel_1956[3];
  assign array_update_1962[4] = sel_1956[4];
  assign array_update_1962[5] = sel_1956[5];
  assign array_update_1962[6] = sgt_1950 ? array_update_1946[add_1898 > 32'h0000_0007 ? 32'h0000_0007 : add_1898] : (sgt_1918 ? array_update_1911[add_1898 > 32'h0000_0007 ? 32'h0000_0007 : add_1898] : (sgt_1881 ? array_update_1875[add_1898 > 32'h0000_0007 ? 32'h0000_0007 : add_1898] : (sgt_1849 ? array_update_1845[add_1898 > 32'h0000_0007 ? 32'h0000_0007 : add_1898] : (sgt_1825 ? array_update_1821[add_1898 > 32'h0000_0007 ? 32'h0000_0007 : add_1898] : (sgt_1804 ? array_update_1803[add_1898 > 32'h0000_0007 ? 32'h0000_0007 : add_1898] : my_string_unflattened[add_1898 > 32'h0000_0007 ? 32'h0000_0007 : add_1898])))));
  assign array_update_1962[7] = sel_1956[7];
  assign array_update_1965[0] = add_1898 == 32'h0000_0000 ? (sgt_1950 ? array_update_1946[3'h6] : (sgt_1918 ? array_update_1911[3'h6] : (sgt_1881 ? array_update_1875[3'h6] : (sgt_1849 ? array_update_1845[3'h6] : (sgt_1825 ? array_update_1821[3'h6] : (sgt_1804 ? array_update_1803[3'h6] : array_index_1736)))))) : array_update_1962[0];
  assign array_update_1965[1] = add_1898 == 32'h0000_0001 ? (sgt_1950 ? array_update_1946[3'h6] : (sgt_1918 ? array_update_1911[3'h6] : (sgt_1881 ? array_update_1875[3'h6] : (sgt_1849 ? array_update_1845[3'h6] : (sgt_1825 ? array_update_1821[3'h6] : (sgt_1804 ? array_update_1803[3'h6] : array_index_1736)))))) : array_update_1962[1];
  assign array_update_1965[2] = add_1898 == 32'h0000_0002 ? (sgt_1950 ? array_update_1946[3'h6] : (sgt_1918 ? array_update_1911[3'h6] : (sgt_1881 ? array_update_1875[3'h6] : (sgt_1849 ? array_update_1845[3'h6] : (sgt_1825 ? array_update_1821[3'h6] : (sgt_1804 ? array_update_1803[3'h6] : array_index_1736)))))) : array_update_1962[2];
  assign array_update_1965[3] = add_1898 == 32'h0000_0003 ? (sgt_1950 ? array_update_1946[3'h6] : (sgt_1918 ? array_update_1911[3'h6] : (sgt_1881 ? array_update_1875[3'h6] : (sgt_1849 ? array_update_1845[3'h6] : (sgt_1825 ? array_update_1821[3'h6] : (sgt_1804 ? array_update_1803[3'h6] : array_index_1736)))))) : array_update_1962[3];
  assign array_update_1965[4] = add_1898 == 32'h0000_0004 ? (sgt_1950 ? array_update_1946[3'h6] : (sgt_1918 ? array_update_1911[3'h6] : (sgt_1881 ? array_update_1875[3'h6] : (sgt_1849 ? array_update_1845[3'h6] : (sgt_1825 ? array_update_1821[3'h6] : (sgt_1804 ? array_update_1803[3'h6] : array_index_1736)))))) : array_update_1962[4];
  assign array_update_1965[5] = add_1898 == 32'h0000_0005 ? (sgt_1950 ? array_update_1946[3'h6] : (sgt_1918 ? array_update_1911[3'h6] : (sgt_1881 ? array_update_1875[3'h6] : (sgt_1849 ? array_update_1845[3'h6] : (sgt_1825 ? array_update_1821[3'h6] : (sgt_1804 ? array_update_1803[3'h6] : array_index_1736)))))) : array_update_1962[5];
  assign array_update_1965[6] = add_1898 == 32'h0000_0006 ? (sgt_1950 ? array_update_1946[3'h6] : (sgt_1918 ? array_update_1911[3'h6] : (sgt_1881 ? array_update_1875[3'h6] : (sgt_1849 ? array_update_1845[3'h6] : (sgt_1825 ? array_update_1821[3'h6] : (sgt_1804 ? array_update_1803[3'h6] : array_index_1736)))))) : array_update_1962[6];
  assign array_update_1965[7] = add_1898 == 32'h0000_0007 ? (sgt_1950 ? array_update_1946[3'h6] : (sgt_1918 ? array_update_1911[3'h6] : (sgt_1881 ? array_update_1875[3'h6] : (sgt_1849 ? array_update_1845[3'h6] : (sgt_1825 ? array_update_1821[3'h6] : (sgt_1804 ? array_update_1803[3'h6] : array_index_1736)))))) : array_update_1962[7];
  assign sel_1966[0] = $signed(and_1790[4:1]) > $signed(4'h6) == 1'h0 ? sel_1956[0] : array_update_1965[0];
  assign sel_1966[1] = $signed(and_1790[4:1]) > $signed(4'h6) == 1'h0 ? sel_1956[1] : array_update_1965[1];
  assign sel_1966[2] = $signed(and_1790[4:1]) > $signed(4'h6) == 1'h0 ? sel_1956[2] : array_update_1965[2];
  assign sel_1966[3] = $signed(and_1790[4:1]) > $signed(4'h6) == 1'h0 ? sel_1956[3] : array_update_1965[3];
  assign sel_1966[4] = $signed(and_1790[4:1]) > $signed(4'h6) == 1'h0 ? sel_1956[4] : array_update_1965[4];
  assign sel_1966[5] = $signed(and_1790[4:1]) > $signed(4'h6) == 1'h0 ? sel_1956[5] : array_update_1965[5];
  assign sel_1966[6] = $signed(and_1790[4:1]) > $signed(4'h6) == 1'h0 ? sel_1956[6] : array_update_1965[6];
  assign sel_1966[7] = $signed(and_1790[4:1]) > $signed(4'h6) == 1'h0 ? sel_1956[7] : array_update_1965[7];
  assign out = {sel_1966[7], sel_1966[6], sel_1966[5], sel_1966[4], sel_1966[3], sel_1966[2], sel_1966[1], sel_1966[0]};
endmodule
